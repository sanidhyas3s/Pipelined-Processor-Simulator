module Program_Counter();
    integer PC;
    initial PC=0;
endmodule