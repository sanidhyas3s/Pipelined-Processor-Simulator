module jump_stall();
    integer js;
    initial js=0;
endmodule