module Memory();
    integer Data[1023:0];
endmodule